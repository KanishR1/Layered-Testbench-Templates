package mac_tb_pkg;

  `include "defines.svh"
  `include "transaction.sv"
  `include "generator.sv"
  `include "driver.sv"
  `include "monitor.sv"
  `include "scoreboard.sv"
  `include "environment.sv"
endpackage