`define DWIDTH 16